module adder_n (input [64:0] a, input [64:0] b, input cin, output [64:0] sum, output cout);
    wire [64:0] carry;

    adder FA0 (a[0], b[0], cin, sum[0], carry[0]);
    adder FA1 (a[1], b[1], carry[0], sum[1], carry[1]);
    adder FA2 (a[2], b[2], carry[1], sum[2], carry[2]);
    adder FA3 (a[3], b[3], carry[2], sum[3], carry[3]);
    adder FA4 (a[4], b[4], carry[3], sum[4], carry[4]);
    adder FA5 (a[5], b[5], carry[4], sum[5], carry[5]);
    adder FA6 (a[6], b[6], carry[5], sum[6], carry[6]);
    adder FA7 (a[7], b[7], carry[6], sum[7], carry[7]);
    adder FA8 (a[8], b[8], carry[7], sum[8], carry[8]);
    adder FA9 (a[9], b[9], carry[8], sum[9], carry[9]);
    adder FA10 (a[10], b[10], carry[9], sum[10], carry[10]);
    adder FA11 (a[11], b[11], carry[10], sum[11], carry[11]);
    adder FA12 (a[12], b[12], carry[11], sum[12], carry[12]);
    adder FA13 (a[13], b[13], carry[12], sum[13], carry[13]);
    adder FA14 (a[14], b[14], carry[13], sum[14], carry[14]);
    adder FA15 (a[15], b[15], carry[14], sum[15], carry[15]);
    adder FA16 (a[16], b[16], carry[15], sum[16], carry[16]);
    adder FA17 (a[17], b[17], carry[16], sum[17], carry[17]);
    adder FA18 (a[18], b[18], carry[17], sum[18], carry[18]);
    adder FA19 (a[19], b[19], carry[18], sum[19], carry[19]);
    adder FA20 (a[20], b[20], carry[19], sum[20], carry[20]);
    adder FA21 (a[21], b[21], carry[20], sum[21], carry[21]);
    adder FA22 (a[22], b[22], carry[21], sum[22], carry[22]);
    adder FA23 (a[23], b[23], carry[22], sum[23], carry[23]);
    adder FA24 (a[24], b[24], carry[23], sum[24], carry[24]);
    adder FA25 (a[25], b[25], carry[24], sum[25], carry[25]);
    adder FA26 (a[26], b[26], carry[25], sum[26], carry[26]);
    adder FA27 (a[27], b[27], carry[26], sum[27], carry[27]);
    adder FA28 (a[28], b[28], carry[27], sum[28], carry[28]);
    adder FA29 (a[29], b[29], carry[28], sum[29], carry[29]);
    adder FA30 (a[30], b[30], carry[29], sum[30], carry[30]);
    adder FA31 (a[31], b[31], carry[30], sum[31], carry[31]);
    adder FA32 (a[32], b[32], carry[31], sum[32], carry[32]);
    adder FA33 (a[33], b[33], carry[32], sum[33], carry[33]);
    adder FA34 (a[34], b[34], carry[33], sum[34], carry[34]);
    adder FA35 (a[35], b[35], carry[34], sum[35], carry[35]);
    adder FA36 (a[36], b[36], carry[35], sum[36], carry[36]);
    adder FA37 (a[37], b[37], carry[36], sum[37], carry[37]);
    adder FA38 (a[38], b[38], carry[37], sum[38], carry[38]);
    adder FA39 (a[39], b[39], carry[38], sum[39], carry[39]);
    adder FA40 (a[40], b[40], carry[39], sum[40], carry[40]);
    adder FA41 (a[41], b[41], carry[40], sum[41], carry[41]);
    adder FA42 (a[42], b[42], carry[41], sum[42], carry[42]);
    adder FA43 (a[43], b[43], carry[42], sum[43], carry[43]);
    adder FA44 (a[44], b[44], carry[43], sum[44], carry[44]);
    adder FA45 (a[45], b[45], carry[44], sum[45], carry[45]);
    adder FA46 (a[46], b[46], carry[45], sum[46], carry[46]);
    adder FA47 (a[47], b[47], carry[46], sum[47], carry[47]);
    adder FA48 (a[48], b[48], carry[47], sum[48], carry[48]);
    adder FA49 (a[49], b[49], carry[48], sum[49], carry[49]);
    adder FA50 (a[50], b[50], carry[49], sum[50], carry[50]);
    adder FA51 (a[51], b[51], carry[50], sum[51], carry[51]);
    adder FA52 (a[52], b[52], carry[51], sum[52], carry[52]);
    adder FA53 (a[53], b[53], carry[52], sum[53], carry[53]);
    adder FA54 (a[54], b[54], carry[53], sum[54], carry[54]);
    adder FA55 (a[55], b[55], carry[54], sum[55], carry[55]);
    adder FA56 (a[56], b[56], carry[55], sum[56], carry[56]);
    adder FA57 (a[57], b[57], carry[56], sum[57], carry[57]);
    adder FA58 (a[58], b[58], carry[57], sum[58], carry[58]);
    adder FA59 (a[59], b[59], carry[58], sum[59], carry[59]);
    adder FA60 (a[60], b[60], carry[59], sum[60], carry[60]);
    adder FA61 (a[61], b[61], carry[60], sum[61], carry[61]);
    adder FA62 (a[62], b[62], carry[61], sum[62], carry[62]);
    adder FA63 (a[63], b[63], carry[62], sum[63], cout);
endmodule